package router_test_pkg;

  int run_for_n_packets = 0;
  int TRACE_ON = 0; 
  `include "router_test.svh"
  `include "Packet.sv"
  `include "Driver.sv"
  `include "Receiver.sv"
  `include "Generator.sv"
  `include "Scoreboard.sv"
  `include "Environment.sv"

endpackage: router_test_pkg