typedef class Packet; // forward typedef
typedef mailbox #(Packet) pkt_mbox;